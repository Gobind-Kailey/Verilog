


module top_module
(
    input wire clk,
    input wire areset,
    input wire in,
    
    
    output reg out
); 

reg [1:0] state, next_state; 

parameter A = 2'b00, B = 2'b01, C = 2'b10, D = 2'b11; 

always@(posedge clk or posedge areset) begin 

    if(areset) state <= A; 
    else state <= next_state; 

end 

always@(*) begin 

    case(state)

 A : next_state = (in)? B : A; 
 B : next_state = (in)? B : C; 
 C : next_state = (in)? D : A; 
 D : next_state = (in)? B : C; 
 default: next_state <= A; 

    endcase

end 
always@(*) begin 

    out = (state == D); 

end 


endmodule