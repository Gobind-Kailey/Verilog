

// We have 2 states: IDLE and Active 
// We an input which is called "start" 
    // When = 1, it will go to active state, otherwise IDLE


module fsm_2_state(
    // State inputs and outputs 

    
    input wire clk, 
    input wire rst, 
    output reg [1:0]
    

)





endmodule