


/*




*/


module top_module
(
    input wire[1:0] state,
    input 
    input wire in,
    output reg q, 



);


endmodule 