



/*

Write Verilog to swap the contents of two registers without using a temporary 
register (and also with a temporary). Then explain how these differ in synthesizable 
logic.

*/


module swap
(

    

);

endmodule 